 -------------------------------------------------------------------------------
-- Copyright (C) 2009 OutputLogic.com
-- This source file may be used and distributed without restriction
-- provided that this copyright statement is not removed from the file
-- and that any derivative work contains the original copyright notice
-- and the associated disclaimer.
--
-- THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
-- WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pkg_hash is
	function hash(slv : std_ulogic_vector) return std_ulogic_vector;
end;

package body pkg_hash is
	function hash(slv : std_ulogic_vector) return std_ulogic_vector is
		variable ret : std_ulogic_vector(11 downto 0) := (others => '1');
	begin
		if slv'length = 296 then
			-- 1 + x^1 + x^3 +x^11 + x^12;
			ret(0)  := slv(0) xor slv(1) xor slv(2) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(10) xor slv(11) xor slv(13) xor slv(15) xor slv(17) xor slv(18) xor slv(21) xor slv(23) xor slv(24) xor slv(28) xor slv(29) xor slv(30) xor slv(31) xor slv(32) xor slv(33) xor slv(36) xor slv(38) xor slv(39) xor slv(41) xor slv(49) xor slv(51) xor slv(53) xor slv(54) xor slv(55) xor slv(56) xor slv(57) xor slv(61) xor slv(62) xor slv(63) xor slv(64) xor slv(66) xor slv(67) xor slv(68) xor slv(70) xor slv(73) xor slv(74) xor slv(79) xor slv(81) xor slv(82) xor slv(84) xor slv(85) xor slv(88) xor slv(89) xor slv(90) xor slv(91) xor slv(93) xor slv(94) xor slv(98) xor slv(99) xor slv(102) xor slv(103) xor slv(106) xor slv(108) xor slv(112) xor slv(118) xor slv(120) xor slv(123) xor slv(127) xor slv(128) xor slv(129) xor slv(131) xor slv(132) xor slv(133) xor slv(135) xor slv(137) xor slv(138) xor slv(139) xor slv(144) xor slv(151) xor slv(152) xor slv(155) xor slv(160) xor slv(162) xor slv(163) xor slv(164) xor slv(165) xor slv(167) xor slv(168) xor slv(174) xor slv(175) xor slv(178) xor slv(179) xor slv(183) xor slv(185) xor slv(186) xor slv(187) xor slv(189) xor slv(190) xor slv(192) xor slv(193) xor slv(194) xor slv(195) xor slv(196) xor slv(197) xor slv(200) xor slv(204) xor slv(206) xor slv(207) xor slv(208) xor slv(209) xor slv(210) xor slv(212) xor slv(218) xor slv(221) xor slv(223) xor slv(227) xor slv(228) xor slv(233) xor slv(235) xor slv(237) xor slv(240) xor slv(241) xor slv(245) xor slv(246) xor slv(248) xor slv(249) xor slv(251) xor slv(252) xor slv(254) xor slv(256) xor slv(259) xor slv(262) xor slv(264) xor slv(265) xor slv(267) xor slv(268) xor slv(269) xor slv(275) xor slv(281) xor slv(282) xor slv(283) xor slv(286) xor slv(290);
			ret(1)  := slv(0) xor slv(9) xor slv(10) xor slv(12) xor slv(13) xor slv(14) xor slv(15) xor slv(16) xor slv(17) xor slv(19) xor slv(21) xor slv(22) xor slv(23) xor slv(25) xor slv(28) xor slv(34) xor slv(36) xor slv(37) xor slv(38) xor slv(40) xor slv(41) xor slv(42) xor slv(49) xor slv(50) xor slv(51) xor slv(52) xor slv(53) xor slv(58) xor slv(61) xor slv(65) xor slv(66) xor slv(69) xor slv(70) xor slv(71) xor slv(73) xor slv(75) xor slv(79) xor slv(80) xor slv(81) xor slv(83) xor slv(84) xor slv(86) xor slv(88) xor slv(92) xor slv(93) xor slv(95) xor slv(98) xor slv(100) xor slv(102) xor slv(104) xor slv(106) xor slv(107) xor slv(108) xor slv(109) xor slv(112) xor slv(113) xor slv(118) xor slv(119) xor slv(120) xor slv(121) xor slv(123) xor slv(124) xor slv(127) xor slv(130) xor slv(131) xor slv(134) xor slv(135) xor slv(136) xor slv(137) xor slv(140) xor slv(144) xor slv(145) xor slv(151) xor slv(153) xor slv(155) xor slv(156) xor slv(160) xor slv(161) xor slv(162) xor slv(166) xor slv(167) xor slv(169) xor slv(174) xor slv(176) xor slv(178) xor slv(180) xor slv(183) xor slv(184) xor slv(185) xor slv(188) xor slv(189) xor slv(191) xor slv(192) xor slv(198) xor slv(200) xor slv(201) xor slv(204) xor slv(205) xor slv(206) xor slv(211) xor slv(212) xor slv(213) xor slv(218) xor slv(219) xor slv(221) xor slv(222) xor slv(223) xor slv(224) xor slv(227) xor slv(229) xor slv(233) xor slv(234) xor slv(235) xor slv(236) xor slv(237) xor slv(238) xor slv(240) xor slv(242) xor slv(245) xor slv(247) xor slv(248) xor slv(250) xor slv(251) xor slv(253) xor slv(254) xor slv(255) xor slv(256) xor slv(257) xor slv(259) xor slv(260) xor slv(262) xor slv(263) xor slv(264) xor slv(266) xor slv(267) xor slv(270) xor slv(275) xor slv(276) xor slv(281) xor slv(284) xor slv(286) xor slv(287) xor slv(290) xor slv(291);
			ret(2)  := slv(1) xor slv(10) xor slv(11) xor slv(13) xor slv(14) xor slv(15) xor slv(16) xor slv(17) xor slv(18) xor slv(20) xor slv(22) xor slv(23) xor slv(24) xor slv(26) xor slv(29) xor slv(35) xor slv(37) xor slv(38) xor slv(39) xor slv(41) xor slv(42) xor slv(43) xor slv(50) xor slv(51) xor slv(52) xor slv(53) xor slv(54) xor slv(59) xor slv(62) xor slv(66) xor slv(67) xor slv(70) xor slv(71) xor slv(72) xor slv(74) xor slv(76) xor slv(80) xor slv(81) xor slv(82) xor slv(84) xor slv(85) xor slv(87) xor slv(89) xor slv(93) xor slv(94) xor slv(96) xor slv(99) xor slv(101) xor slv(103) xor slv(105) xor slv(107) xor slv(108) xor slv(109) xor slv(110) xor slv(113) xor slv(114) xor slv(119) xor slv(120) xor slv(121) xor slv(122) xor slv(124) xor slv(125) xor slv(128) xor slv(131) xor slv(132) xor slv(135) xor slv(136) xor slv(137) xor slv(138) xor slv(141) xor slv(145) xor slv(146) xor slv(152) xor slv(154) xor slv(156) xor slv(157) xor slv(161) xor slv(162) xor slv(163) xor slv(167) xor slv(168) xor slv(170) xor slv(175) xor slv(177) xor slv(179) xor slv(181) xor slv(184) xor slv(185) xor slv(186) xor slv(189) xor slv(190) xor slv(192) xor slv(193) xor slv(199) xor slv(201) xor slv(202) xor slv(205) xor slv(206) xor slv(207) xor slv(212) xor slv(213) xor slv(214) xor slv(219) xor slv(220) xor slv(222) xor slv(223) xor slv(224) xor slv(225) xor slv(228) xor slv(230) xor slv(234) xor slv(235) xor slv(236) xor slv(237) xor slv(238) xor slv(239) xor slv(241) xor slv(243) xor slv(246) xor slv(248) xor slv(249) xor slv(251) xor slv(252) xor slv(254) xor slv(255) xor slv(256) xor slv(257) xor slv(258) xor slv(260) xor slv(261) xor slv(263) xor slv(264) xor slv(265) xor slv(267) xor slv(268) xor slv(271) xor slv(276) xor slv(277) xor slv(282) xor slv(285) xor slv(287) xor slv(288) xor slv(291) xor slv(292);
			ret(3)  := slv(0) xor slv(1) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(10) xor slv(12) xor slv(13) xor slv(14) xor slv(16) xor slv(19) xor slv(25) xor slv(27) xor slv(28) xor slv(29) xor slv(31) xor slv(32) xor slv(33) xor slv(40) xor slv(41) xor slv(42) xor slv(43) xor slv(44) xor slv(49) xor slv(52) xor slv(56) xor slv(57) xor slv(60) xor slv(61) xor slv(62) xor slv(64) xor slv(66) xor slv(70) xor slv(71) xor slv(72) xor slv(74) xor slv(75) xor slv(77) xor slv(79) xor slv(83) xor slv(84) xor slv(86) xor slv(89) xor slv(91) xor slv(93) xor slv(95) xor slv(97) xor slv(98) xor slv(99) xor slv(100) xor slv(103) xor slv(104) xor slv(109) xor slv(110) xor slv(111) xor slv(112) xor slv(114) xor slv(115) xor slv(118) xor slv(121) xor slv(122) xor slv(125) xor slv(126) xor slv(127) xor slv(128) xor slv(131) xor slv(135) xor slv(136) xor slv(142) xor slv(144) xor slv(146) xor slv(147) xor slv(151) xor slv(152) xor slv(153) xor slv(157) xor slv(158) xor slv(160) xor slv(165) xor slv(167) xor slv(169) xor slv(171) xor slv(174) xor slv(175) xor slv(176) xor slv(179) xor slv(180) xor slv(182) xor slv(183) xor slv(189) xor slv(191) xor slv(192) xor slv(195) xor slv(196) xor slv(197) xor slv(202) xor slv(203) xor slv(204) xor slv(209) xor slv(210) xor slv(212) xor slv(213) xor slv(214) xor slv(215) xor slv(218) xor slv(220) xor slv(224) xor slv(225) xor slv(226) xor slv(227) xor slv(228) xor slv(229) xor slv(231) xor slv(233) xor slv(236) xor slv(238) xor slv(239) xor slv(241) xor slv(242) xor slv(244) xor slv(245) xor slv(246) xor slv(247) xor slv(248) xor slv(250) xor slv(251) xor slv(253) xor slv(254) xor slv(255) xor slv(257) xor slv(258) xor slv(261) xor slv(266) xor slv(267) xor slv(272) xor slv(275) xor slv(277) xor slv(278) xor slv(281) xor slv(282) xor slv(288) xor slv(289) xor slv(290) xor slv(292) xor slv(293);
			ret(4)  := slv(1) xor slv(2) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(11) xor slv(13) xor slv(14) xor slv(15) xor slv(17) xor slv(20) xor slv(26) xor slv(28) xor slv(29) xor slv(30) xor slv(32) xor slv(33) xor slv(34) xor slv(41) xor slv(42) xor slv(43) xor slv(44) xor slv(45) xor slv(50) xor slv(53) xor slv(57) xor slv(58) xor slv(61) xor slv(62) xor slv(63) xor slv(65) xor slv(67) xor slv(71) xor slv(72) xor slv(73) xor slv(75) xor slv(76) xor slv(78) xor slv(80) xor slv(84) xor slv(85) xor slv(87) xor slv(90) xor slv(92) xor slv(94) xor slv(96) xor slv(98) xor slv(99) xor slv(100) xor slv(101) xor slv(104) xor slv(105) xor slv(110) xor slv(111) xor slv(112) xor slv(113) xor slv(115) xor slv(116) xor slv(119) xor slv(122) xor slv(123) xor slv(126) xor slv(127) xor slv(128) xor slv(129) xor slv(132) xor slv(136) xor slv(137) xor slv(143) xor slv(145) xor slv(147) xor slv(148) xor slv(152) xor slv(153) xor slv(154) xor slv(158) xor slv(159) xor slv(161) xor slv(166) xor slv(168) xor slv(170) xor slv(172) xor slv(175) xor slv(176) xor slv(177) xor slv(180) xor slv(181) xor slv(183) xor slv(184) xor slv(190) xor slv(192) xor slv(193) xor slv(196) xor slv(197) xor slv(198) xor slv(203) xor slv(204) xor slv(205) xor slv(210) xor slv(211) xor slv(213) xor slv(214) xor slv(215) xor slv(216) xor slv(219) xor slv(221) xor slv(225) xor slv(226) xor slv(227) xor slv(228) xor slv(229) xor slv(230) xor slv(232) xor slv(234) xor slv(237) xor slv(239) xor slv(240) xor slv(242) xor slv(243) xor slv(245) xor slv(246) xor slv(247) xor slv(248) xor slv(249) xor slv(251) xor slv(252) xor slv(254) xor slv(255) xor slv(256) xor slv(258) xor slv(259) xor slv(262) xor slv(267) xor slv(268) xor slv(273) xor slv(276) xor slv(278) xor slv(279) xor slv(282) xor slv(283) xor slv(289) xor slv(290) xor slv(291) xor slv(293) xor slv(294);
			ret(5)  := slv(2) xor slv(3) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(12) xor slv(14) xor slv(15) xor slv(16) xor slv(18) xor slv(21) xor slv(27) xor slv(29) xor slv(30) xor slv(31) xor slv(33) xor slv(34) xor slv(35) xor slv(42) xor slv(43) xor slv(44) xor slv(45) xor slv(46) xor slv(51) xor slv(54) xor slv(58) xor slv(59) xor slv(62) xor slv(63) xor slv(64) xor slv(66) xor slv(68) xor slv(72) xor slv(73) xor slv(74) xor slv(76) xor slv(77) xor slv(79) xor slv(81) xor slv(85) xor slv(86) xor slv(88) xor slv(91) xor slv(93) xor slv(95) xor slv(97) xor slv(99) xor slv(100) xor slv(101) xor slv(102) xor slv(105) xor slv(106) xor slv(111) xor slv(112) xor slv(113) xor slv(114) xor slv(116) xor slv(117) xor slv(120) xor slv(123) xor slv(124) xor slv(127) xor slv(128) xor slv(129) xor slv(130) xor slv(133) xor slv(137) xor slv(138) xor slv(144) xor slv(146) xor slv(148) xor slv(149) xor slv(153) xor slv(154) xor slv(155) xor slv(159) xor slv(160) xor slv(162) xor slv(167) xor slv(169) xor slv(171) xor slv(173) xor slv(176) xor slv(177) xor slv(178) xor slv(181) xor slv(182) xor slv(184) xor slv(185) xor slv(191) xor slv(193) xor slv(194) xor slv(197) xor slv(198) xor slv(199) xor slv(204) xor slv(205) xor slv(206) xor slv(211) xor slv(212) xor slv(214) xor slv(215) xor slv(216) xor slv(217) xor slv(220) xor slv(222) xor slv(226) xor slv(227) xor slv(228) xor slv(229) xor slv(230) xor slv(231) xor slv(233) xor slv(235) xor slv(238) xor slv(240) xor slv(241) xor slv(243) xor slv(244) xor slv(246) xor slv(247) xor slv(248) xor slv(249) xor slv(250) xor slv(252) xor slv(253) xor slv(255) xor slv(256) xor slv(257) xor slv(259) xor slv(260) xor slv(263) xor slv(268) xor slv(269) xor slv(274) xor slv(277) xor slv(279) xor slv(280) xor slv(283) xor slv(284) xor slv(290) xor slv(291) xor slv(292) xor slv(294) xor slv(295);
			ret(6)  := slv(3) xor slv(4) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(13) xor slv(15) xor slv(16) xor slv(17) xor slv(19) xor slv(22) xor slv(28) xor slv(30) xor slv(31) xor slv(32) xor slv(34) xor slv(35) xor slv(36) xor slv(43) xor slv(44) xor slv(45) xor slv(46) xor slv(47) xor slv(52) xor slv(55) xor slv(59) xor slv(60) xor slv(63) xor slv(64) xor slv(65) xor slv(67) xor slv(69) xor slv(73) xor slv(74) xor slv(75) xor slv(77) xor slv(78) xor slv(80) xor slv(82) xor slv(86) xor slv(87) xor slv(89) xor slv(92) xor slv(94) xor slv(96) xor slv(98) xor slv(100) xor slv(101) xor slv(102) xor slv(103) xor slv(106) xor slv(107) xor slv(112) xor slv(113) xor slv(114) xor slv(115) xor slv(117) xor slv(118) xor slv(121) xor slv(124) xor slv(125) xor slv(128) xor slv(129) xor slv(130) xor slv(131) xor slv(134) xor slv(138) xor slv(139) xor slv(145) xor slv(147) xor slv(149) xor slv(150) xor slv(154) xor slv(155) xor slv(156) xor slv(160) xor slv(161) xor slv(163) xor slv(168) xor slv(170) xor slv(172) xor slv(174) xor slv(177) xor slv(178) xor slv(179) xor slv(182) xor slv(183) xor slv(185) xor slv(186) xor slv(192) xor slv(194) xor slv(195) xor slv(198) xor slv(199) xor slv(200) xor slv(205) xor slv(206) xor slv(207) xor slv(212) xor slv(213) xor slv(215) xor slv(216) xor slv(217) xor slv(218) xor slv(221) xor slv(223) xor slv(227) xor slv(228) xor slv(229) xor slv(230) xor slv(231) xor slv(232) xor slv(234) xor slv(236) xor slv(239) xor slv(241) xor slv(242) xor slv(244) xor slv(245) xor slv(247) xor slv(248) xor slv(249) xor slv(250) xor slv(251) xor slv(253) xor slv(254) xor slv(256) xor slv(257) xor slv(258) xor slv(260) xor slv(261) xor slv(264) xor slv(269) xor slv(270) xor slv(275) xor slv(278) xor slv(280) xor slv(281) xor slv(284) xor slv(285) xor slv(291) xor slv(292) xor slv(293) xor slv(295);
			ret(7)  := slv(4) xor slv(5) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(14) xor slv(16) xor slv(17) xor slv(18) xor slv(20) xor slv(23) xor slv(29) xor slv(31) xor slv(32) xor slv(33) xor slv(35) xor slv(36) xor slv(37) xor slv(44) xor slv(45) xor slv(46) xor slv(47) xor slv(48) xor slv(53) xor slv(56) xor slv(60) xor slv(61) xor slv(64) xor slv(65) xor slv(66) xor slv(68) xor slv(70) xor slv(74) xor slv(75) xor slv(76) xor slv(78) xor slv(79) xor slv(81) xor slv(83) xor slv(87) xor slv(88) xor slv(90) xor slv(93) xor slv(95) xor slv(97) xor slv(99) xor slv(101) xor slv(102) xor slv(103) xor slv(104) xor slv(107) xor slv(108) xor slv(113) xor slv(114) xor slv(115) xor slv(116) xor slv(118) xor slv(119) xor slv(122) xor slv(125) xor slv(126) xor slv(129) xor slv(130) xor slv(131) xor slv(132) xor slv(135) xor slv(139) xor slv(140) xor slv(146) xor slv(148) xor slv(150) xor slv(151) xor slv(155) xor slv(156) xor slv(157) xor slv(161) xor slv(162) xor slv(164) xor slv(169) xor slv(171) xor slv(173) xor slv(175) xor slv(178) xor slv(179) xor slv(180) xor slv(183) xor slv(184) xor slv(186) xor slv(187) xor slv(193) xor slv(195) xor slv(196) xor slv(199) xor slv(200) xor slv(201) xor slv(206) xor slv(207) xor slv(208) xor slv(213) xor slv(214) xor slv(216) xor slv(217) xor slv(218) xor slv(219) xor slv(222) xor slv(224) xor slv(228) xor slv(229) xor slv(230) xor slv(231) xor slv(232) xor slv(233) xor slv(235) xor slv(237) xor slv(240) xor slv(242) xor slv(243) xor slv(245) xor slv(246) xor slv(248) xor slv(249) xor slv(250) xor slv(251) xor slv(252) xor slv(254) xor slv(255) xor slv(257) xor slv(258) xor slv(259) xor slv(261) xor slv(262) xor slv(265) xor slv(270) xor slv(271) xor slv(276) xor slv(279) xor slv(281) xor slv(282) xor slv(285) xor slv(286) xor slv(292) xor slv(293) xor slv(294);
			ret(8)  := slv(5) xor slv(6) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(15) xor slv(17) xor slv(18) xor slv(19) xor slv(21) xor slv(24) xor slv(30) xor slv(32) xor slv(33) xor slv(34) xor slv(36) xor slv(37) xor slv(38) xor slv(45) xor slv(46) xor slv(47) xor slv(48) xor slv(49) xor slv(54) xor slv(57) xor slv(61) xor slv(62) xor slv(65) xor slv(66) xor slv(67) xor slv(69) xor slv(71) xor slv(75) xor slv(76) xor slv(77) xor slv(79) xor slv(80) xor slv(82) xor slv(84) xor slv(88) xor slv(89) xor slv(91) xor slv(94) xor slv(96) xor slv(98) xor slv(100) xor slv(102) xor slv(103) xor slv(104) xor slv(105) xor slv(108) xor slv(109) xor slv(114) xor slv(115) xor slv(116) xor slv(117) xor slv(119) xor slv(120) xor slv(123) xor slv(126) xor slv(127) xor slv(130) xor slv(131) xor slv(132) xor slv(133) xor slv(136) xor slv(140) xor slv(141) xor slv(147) xor slv(149) xor slv(151) xor slv(152) xor slv(156) xor slv(157) xor slv(158) xor slv(162) xor slv(163) xor slv(165) xor slv(170) xor slv(172) xor slv(174) xor slv(176) xor slv(179) xor slv(180) xor slv(181) xor slv(184) xor slv(185) xor slv(187) xor slv(188) xor slv(194) xor slv(196) xor slv(197) xor slv(200) xor slv(201) xor slv(202) xor slv(207) xor slv(208) xor slv(209) xor slv(214) xor slv(215) xor slv(217) xor slv(218) xor slv(219) xor slv(220) xor slv(223) xor slv(225) xor slv(229) xor slv(230) xor slv(231) xor slv(232) xor slv(233) xor slv(234) xor slv(236) xor slv(238) xor slv(241) xor slv(243) xor slv(244) xor slv(246) xor slv(247) xor slv(249) xor slv(250) xor slv(251) xor slv(252) xor slv(253) xor slv(255) xor slv(256) xor slv(258) xor slv(259) xor slv(260) xor slv(262) xor slv(263) xor slv(266) xor slv(271) xor slv(272) xor slv(277) xor slv(280) xor slv(282) xor slv(283) xor slv(286) xor slv(287) xor slv(293) xor slv(294) xor slv(295);
			ret(9)  := slv(6) xor slv(7) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(14) xor slv(16) xor slv(18) xor slv(19) xor slv(20) xor slv(22) xor slv(25) xor slv(31) xor slv(33) xor slv(34) xor slv(35) xor slv(37) xor slv(38) xor slv(39) xor slv(46) xor slv(47) xor slv(48) xor slv(49) xor slv(50) xor slv(55) xor slv(58) xor slv(62) xor slv(63) xor slv(66) xor slv(67) xor slv(68) xor slv(70) xor slv(72) xor slv(76) xor slv(77) xor slv(78) xor slv(80) xor slv(81) xor slv(83) xor slv(85) xor slv(89) xor slv(90) xor slv(92) xor slv(95) xor slv(97) xor slv(99) xor slv(101) xor slv(103) xor slv(104) xor slv(105) xor slv(106) xor slv(109) xor slv(110) xor slv(115) xor slv(116) xor slv(117) xor slv(118) xor slv(120) xor slv(121) xor slv(124) xor slv(127) xor slv(128) xor slv(131) xor slv(132) xor slv(133) xor slv(134) xor slv(137) xor slv(141) xor slv(142) xor slv(148) xor slv(150) xor slv(152) xor slv(153) xor slv(157) xor slv(158) xor slv(159) xor slv(163) xor slv(164) xor slv(166) xor slv(171) xor slv(173) xor slv(175) xor slv(177) xor slv(180) xor slv(181) xor slv(182) xor slv(185) xor slv(186) xor slv(188) xor slv(189) xor slv(195) xor slv(197) xor slv(198) xor slv(201) xor slv(202) xor slv(203) xor slv(208) xor slv(209) xor slv(210) xor slv(215) xor slv(216) xor slv(218) xor slv(219) xor slv(220) xor slv(221) xor slv(224) xor slv(226) xor slv(230) xor slv(231) xor slv(232) xor slv(233) xor slv(234) xor slv(235) xor slv(237) xor slv(239) xor slv(242) xor slv(244) xor slv(245) xor slv(247) xor slv(248) xor slv(250) xor slv(251) xor slv(252) xor slv(253) xor slv(254) xor slv(256) xor slv(257) xor slv(259) xor slv(260) xor slv(261) xor slv(263) xor slv(264) xor slv(267) xor slv(272) xor slv(273) xor slv(278) xor slv(281) xor slv(283) xor slv(284) xor slv(287) xor slv(288) xor slv(294) xor slv(295);
			ret(10) := slv(7) xor slv(8) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(14) xor slv(15) xor slv(17) xor slv(19) xor slv(20) xor slv(21) xor slv(23) xor slv(26) xor slv(32) xor slv(34) xor slv(35) xor slv(36) xor slv(38) xor slv(39) xor slv(40) xor slv(47) xor slv(48) xor slv(49) xor slv(50) xor slv(51) xor slv(56) xor slv(59) xor slv(63) xor slv(64) xor slv(67) xor slv(68) xor slv(69) xor slv(71) xor slv(73) xor slv(77) xor slv(78) xor slv(79) xor slv(81) xor slv(82) xor slv(84) xor slv(86) xor slv(90) xor slv(91) xor slv(93) xor slv(96) xor slv(98) xor slv(100) xor slv(102) xor slv(104) xor slv(105) xor slv(106) xor slv(107) xor slv(110) xor slv(111) xor slv(116) xor slv(117) xor slv(118) xor slv(119) xor slv(121) xor slv(122) xor slv(125) xor slv(128) xor slv(129) xor slv(132) xor slv(133) xor slv(134) xor slv(135) xor slv(138) xor slv(142) xor slv(143) xor slv(149) xor slv(151) xor slv(153) xor slv(154) xor slv(158) xor slv(159) xor slv(160) xor slv(164) xor slv(165) xor slv(167) xor slv(172) xor slv(174) xor slv(176) xor slv(178) xor slv(181) xor slv(182) xor slv(183) xor slv(186) xor slv(187) xor slv(189) xor slv(190) xor slv(196) xor slv(198) xor slv(199) xor slv(202) xor slv(203) xor slv(204) xor slv(209) xor slv(210) xor slv(211) xor slv(216) xor slv(217) xor slv(219) xor slv(220) xor slv(221) xor slv(222) xor slv(225) xor slv(227) xor slv(231) xor slv(232) xor slv(233) xor slv(234) xor slv(235) xor slv(236) xor slv(238) xor slv(240) xor slv(243) xor slv(245) xor slv(246) xor slv(248) xor slv(249) xor slv(251) xor slv(252) xor slv(253) xor slv(254) xor slv(255) xor slv(257) xor slv(258) xor slv(260) xor slv(261) xor slv(262) xor slv(264) xor slv(265) xor slv(268) xor slv(273) xor slv(274) xor slv(279) xor slv(282) xor slv(284) xor slv(285) xor slv(288) xor slv(289) xor slv(295);
			ret(11) := slv(0) xor slv(1) xor slv(2) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(9) xor slv(10) xor slv(12) xor slv(14) xor slv(16) xor slv(17) xor slv(20) xor slv(22) xor slv(23) xor slv(27) xor slv(28) xor slv(29) xor slv(30) xor slv(31) xor slv(32) xor slv(35) xor slv(37) xor slv(38) xor slv(40) xor slv(48) xor slv(50) xor slv(52) xor slv(53) xor slv(54) xor slv(55) xor slv(56) xor slv(60) xor slv(61) xor slv(62) xor slv(63) xor slv(65) xor slv(66) xor slv(67) xor slv(69) xor slv(72) xor slv(73) xor slv(78) xor slv(80) xor slv(81) xor slv(83) xor slv(84) xor slv(87) xor slv(88) xor slv(89) xor slv(90) xor slv(92) xor slv(93) xor slv(97) xor slv(98) xor slv(101) xor slv(102) xor slv(105) xor slv(107) xor slv(111) xor slv(117) xor slv(119) xor slv(122) xor slv(126) xor slv(127) xor slv(128) xor slv(130) xor slv(131) xor slv(132) xor slv(134) xor slv(136) xor slv(137) xor slv(138) xor slv(143) xor slv(150) xor slv(151) xor slv(154) xor slv(159) xor slv(161) xor slv(162) xor slv(163) xor slv(164) xor slv(166) xor slv(167) xor slv(173) xor slv(174) xor slv(177) xor slv(178) xor slv(182) xor slv(184) xor slv(185) xor slv(186) xor slv(188) xor slv(189) xor slv(191) xor slv(192) xor slv(193) xor slv(194) xor slv(195) xor slv(196) xor slv(199) xor slv(203) xor slv(205) xor slv(206) xor slv(207) xor slv(208) xor slv(209) xor slv(211) xor slv(217) xor slv(220) xor slv(222) xor slv(226) xor slv(227) xor slv(232) xor slv(234) xor slv(236) xor slv(239) xor slv(240) xor slv(244) xor slv(245) xor slv(247) xor slv(248) xor slv(250) xor slv(251) xor slv(253) xor slv(255) xor slv(258) xor slv(261) xor slv(263) xor slv(264) xor slv(266) xor slv(267) xor slv(268) xor slv(274) xor slv(280) xor slv(281) xor slv(282) xor slv(285) xor slv(289);
			return ret;
		elsif slv'length = 104 then
			-- 1 + x^1 + x^3 + x^11 + x^12;
			ret(0)  := slv(0) xor slv(1) xor slv(2) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(10) xor slv(11) xor slv(13) xor slv(15) xor slv(17) xor slv(18) xor slv(21) xor slv(23) xor slv(24) xor slv(28) xor slv(29) xor slv(30) xor slv(31) xor slv(32) xor slv(33) xor slv(36) xor slv(38) xor slv(39) xor slv(41) xor slv(49) xor slv(51) xor slv(53) xor slv(54) xor slv(55) xor slv(56) xor slv(57) xor slv(61) xor slv(62) xor slv(63) xor slv(64) xor slv(66) xor slv(67) xor slv(68) xor slv(70) xor slv(73) xor slv(74) xor slv(79) xor slv(81) xor slv(82) xor slv(84) xor slv(85) xor slv(88) xor slv(89) xor slv(90) xor slv(91) xor slv(93) xor slv(94) xor slv(98) xor slv(99) xor slv(102) xor slv(103);
			ret(1)  := slv(0) xor slv(9) xor slv(10) xor slv(12) xor slv(13) xor slv(14) xor slv(15) xor slv(16) xor slv(17) xor slv(19) xor slv(21) xor slv(22) xor slv(23) xor slv(25) xor slv(28) xor slv(34) xor slv(36) xor slv(37) xor slv(38) xor slv(40) xor slv(41) xor slv(42) xor slv(49) xor slv(50) xor slv(51) xor slv(52) xor slv(53) xor slv(58) xor slv(61) xor slv(65) xor slv(66) xor slv(69) xor slv(70) xor slv(71) xor slv(73) xor slv(75) xor slv(79) xor slv(80) xor slv(81) xor slv(83) xor slv(84) xor slv(86) xor slv(88) xor slv(92) xor slv(93) xor slv(95) xor slv(98) xor slv(100) xor slv(102);
			ret(2)  := slv(1) xor slv(10) xor slv(11) xor slv(13) xor slv(14) xor slv(15) xor slv(16) xor slv(17) xor slv(18) xor slv(20) xor slv(22) xor slv(23) xor slv(24) xor slv(26) xor slv(29) xor slv(35) xor slv(37) xor slv(38) xor slv(39) xor slv(41) xor slv(42) xor slv(43) xor slv(50) xor slv(51) xor slv(52) xor slv(53) xor slv(54) xor slv(59) xor slv(62) xor slv(66) xor slv(67) xor slv(70) xor slv(71) xor slv(72) xor slv(74) xor slv(76) xor slv(80) xor slv(81) xor slv(82) xor slv(84) xor slv(85) xor slv(87) xor slv(89) xor slv(93) xor slv(94) xor slv(96) xor slv(99) xor slv(101) xor slv(103);
			ret(3)  := slv(0) xor slv(1) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(10) xor slv(12) xor slv(13) xor slv(14) xor slv(16) xor slv(19) xor slv(25) xor slv(27) xor slv(28) xor slv(29) xor slv(31) xor slv(32) xor slv(33) xor slv(40) xor slv(41) xor slv(42) xor slv(43) xor slv(44) xor slv(49) xor slv(52) xor slv(56) xor slv(57) xor slv(60) xor slv(61) xor slv(62) xor slv(64) xor slv(66) xor slv(70) xor slv(71) xor slv(72) xor slv(74) xor slv(75) xor slv(77) xor slv(79) xor slv(83) xor slv(84) xor slv(86) xor slv(89) xor slv(91) xor slv(93) xor slv(95) xor slv(97) xor slv(98) xor slv(99) xor slv(100) xor slv(103);
			ret(4)  := slv(1) xor slv(2) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(11) xor slv(13) xor slv(14) xor slv(15) xor slv(17) xor slv(20) xor slv(26) xor slv(28) xor slv(29) xor slv(30) xor slv(32) xor slv(33) xor slv(34) xor slv(41) xor slv(42) xor slv(43) xor slv(44) xor slv(45) xor slv(50) xor slv(53) xor slv(57) xor slv(58) xor slv(61) xor slv(62) xor slv(63) xor slv(65) xor slv(67) xor slv(71) xor slv(72) xor slv(73) xor slv(75) xor slv(76) xor slv(78) xor slv(80) xor slv(84) xor slv(85) xor slv(87) xor slv(90) xor slv(92) xor slv(94) xor slv(96) xor slv(98) xor slv(99) xor slv(100) xor slv(101);
			ret(5)  := slv(2) xor slv(3) xor slv(5) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(12) xor slv(14) xor slv(15) xor slv(16) xor slv(18) xor slv(21) xor slv(27) xor slv(29) xor slv(30) xor slv(31) xor slv(33) xor slv(34) xor slv(35) xor slv(42) xor slv(43) xor slv(44) xor slv(45) xor slv(46) xor slv(51) xor slv(54) xor slv(58) xor slv(59) xor slv(62) xor slv(63) xor slv(64) xor slv(66) xor slv(68) xor slv(72) xor slv(73) xor slv(74) xor slv(76) xor slv(77) xor slv(79) xor slv(81) xor slv(85) xor slv(86) xor slv(88) xor slv(91) xor slv(93) xor slv(95) xor slv(97) xor slv(99) xor slv(100) xor slv(101) xor slv(102);
			ret(6)  := slv(3) xor slv(4) xor slv(6) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(13) xor slv(15) xor slv(16) xor slv(17) xor slv(19) xor slv(22) xor slv(28) xor slv(30) xor slv(31) xor slv(32) xor slv(34) xor slv(35) xor slv(36) xor slv(43) xor slv(44) xor slv(45) xor slv(46) xor slv(47) xor slv(52) xor slv(55) xor slv(59) xor slv(60) xor slv(63) xor slv(64) xor slv(65) xor slv(67) xor slv(69) xor slv(73) xor slv(74) xor slv(75) xor slv(77) xor slv(78) xor slv(80) xor slv(82) xor slv(86) xor slv(87) xor slv(89) xor slv(92) xor slv(94) xor slv(96) xor slv(98) xor slv(100) xor slv(101) xor slv(102) xor slv(103);
			ret(7)  := slv(4) xor slv(5) xor slv(7) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(14) xor slv(16) xor slv(17) xor slv(18) xor slv(20) xor slv(23) xor slv(29) xor slv(31) xor slv(32) xor slv(33) xor slv(35) xor slv(36) xor slv(37) xor slv(44) xor slv(45) xor slv(46) xor slv(47) xor slv(48) xor slv(53) xor slv(56) xor slv(60) xor slv(61) xor slv(64) xor slv(65) xor slv(66) xor slv(68) xor slv(70) xor slv(74) xor slv(75) xor slv(76) xor slv(78) xor slv(79) xor slv(81) xor slv(83) xor slv(87) xor slv(88) xor slv(90) xor slv(93) xor slv(95) xor slv(97) xor slv(99) xor slv(101) xor slv(102) xor slv(103);
			ret(8)  := slv(5) xor slv(6) xor slv(8) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(15) xor slv(17) xor slv(18) xor slv(19) xor slv(21) xor slv(24) xor slv(30) xor slv(32) xor slv(33) xor slv(34) xor slv(36) xor slv(37) xor slv(38) xor slv(45) xor slv(46) xor slv(47) xor slv(48) xor slv(49) xor slv(54) xor slv(57) xor slv(61) xor slv(62) xor slv(65) xor slv(66) xor slv(67) xor slv(69) xor slv(71) xor slv(75) xor slv(76) xor slv(77) xor slv(79) xor slv(80) xor slv(82) xor slv(84) xor slv(88) xor slv(89) xor slv(91) xor slv(94) xor slv(96) xor slv(98) xor slv(100) xor slv(102) xor slv(103);
			ret(9)  := slv(6) xor slv(7) xor slv(9) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(14) xor slv(16) xor slv(18) xor slv(19) xor slv(20) xor slv(22) xor slv(25) xor slv(31) xor slv(33) xor slv(34) xor slv(35) xor slv(37) xor slv(38) xor slv(39) xor slv(46) xor slv(47) xor slv(48) xor slv(49) xor slv(50) xor slv(55) xor slv(58) xor slv(62) xor slv(63) xor slv(66) xor slv(67) xor slv(68) xor slv(70) xor slv(72) xor slv(76) xor slv(77) xor slv(78) xor slv(80) xor slv(81) xor slv(83) xor slv(85) xor slv(89) xor slv(90) xor slv(92) xor slv(95) xor slv(97) xor slv(99) xor slv(101) xor slv(103);
			ret(10) := slv(7) xor slv(8) xor slv(10) xor slv(11) xor slv(12) xor slv(13) xor slv(14) xor slv(15) xor slv(17) xor slv(19) xor slv(20) xor slv(21) xor slv(23) xor slv(26) xor slv(32) xor slv(34) xor slv(35) xor slv(36) xor slv(38) xor slv(39) xor slv(40) xor slv(47) xor slv(48) xor slv(49) xor slv(50) xor slv(51) xor slv(56) xor slv(59) xor slv(63) xor slv(64) xor slv(67) xor slv(68) xor slv(69) xor slv(71) xor slv(73) xor slv(77) xor slv(78) xor slv(79) xor slv(81) xor slv(82) xor slv(84) xor slv(86) xor slv(90) xor slv(91) xor slv(93) xor slv(96) xor slv(98) xor slv(100) xor slv(102);
			ret(11) := slv(0) xor slv(1) xor slv(2) xor slv(3) xor slv(4) xor slv(5) xor slv(6) xor slv(7) xor slv(9) xor slv(10) xor slv(12) xor slv(14) xor slv(16) xor slv(17) xor slv(20) xor slv(22) xor slv(23) xor slv(27) xor slv(28) xor slv(29) xor slv(30) xor slv(31) xor slv(32) xor slv(35) xor slv(37) xor slv(38) xor slv(40) xor slv(48) xor slv(50) xor slv(52) xor slv(53) xor slv(54) xor slv(55) xor slv(56) xor slv(60) xor slv(61) xor slv(62) xor slv(63) xor slv(65) xor slv(66) xor slv(67) xor slv(69) xor slv(72) xor slv(73) xor slv(78) xor slv(80) xor slv(81) xor slv(83) xor slv(84) xor slv(87) xor slv(88) xor slv(89) xor slv(90) xor slv(92) xor slv(93) xor slv(97) xor slv(98) xor slv(101) xor slv(102);
			return ret;
		else
			assert false
				report "hash function not defined for input width " & integer'image(slv'length)
				severity failure;
			return x"000";
		end if;
	end;
end;
